** sch_path: /foss/designs/unic-cass-dpga/xschem/Ota_cmrr_tb.sch
**.subckt Ota_cmrr_tb
x1 net1 in ip out net2 GND Ota_esq
Vip ip GND DC 0.9 AC 1
.save i(vip)
VDD net1 GND 1.8
.save i(vdd)
I0 net2 GND 15u
x2 net3 cmrr cmrr out2 net4 GND Ota_esq
Vcmrr cmrr GND DC 0.9 AC 1
.save i(vcmrr)
VDD2 net3 GND 1.8
.save i(vdd2)
I1 net4 GND 15u
Vin in GND DC 0.9 AC 1 180
.save i(vin)
C1 out GND 4p m=1
C2 out2 GND 4p m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt



*cmd step stop

.ac dec 2000 1 110Meg
.save all
.end

.control
run
*CMRR
let cmrr = db((v(out)/(v(ip)-v(in)))/(v(out2)/v(cmrr)))
plot cmrr
*plot db((v(out)/(v(ip)-v(in)))/(v(out2)/v(cmrr)))
*Ganho de modo comum
let mod_com = db(v(out2)/v(cmrr))
plot mod_com
*plot db(v(out2)/v(cmrr))
*Ganho diferencial
let mod_dif = db(v(out)/(v(ip)-v(in)))
plot mod_dif
*plot db(v(out)/(v(ip)-v(in)))
.endc

**** end user architecture code
**.ends

* expanding   symbol:  Ota_esq.sym # of pins=6
** sym_path: /foss/designs/unic-cass-dpga/xschem/Ota_esq.sym
** sch_path: /foss/designs/unic-cass-dpga/xschem/Ota_esq.sch
.subckt Ota_esq VDD Vin Vip Vout Ibias VSS
*.ipin Vin
*.ipin Vip
*.iopin VDD
*.iopin VSS
*.iopin Ibias
*.opin Vout
XM1 net1 Vin net3 net3 sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 Vip net3 net3 sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=8 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=8 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net3 Ibias VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=24 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 Ibias Ibias VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=24 nf=8 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vout Ibias VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=39 nf=13 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout net2 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=21 nf=7 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC1 net2 Vout sky130_fd_pr__cap_mim_m3_1 W=23 L=23 MF=1 m=1
.ends

.GLOBAL GND
.end
